////ody shbayeh left shift reg//// 
////project_1201462////

module leftshift_ody_1201462 #(parameter n=3) (x,y);///module 
input signed [n:0] x ;///input
output reg signed [n+1:0] y ;//output

always @(x) ///shift left by 1 bit as a multiplication by 2
 begin 
 
 y = x*2;
 end 
 
 endmodule 